module rr_arb
(
  input clk,
)

endmodule
